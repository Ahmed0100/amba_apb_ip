`define IP_AMBA_APB_MASTER_PARAM_DECL #(parameter PRDATA_width = `PRDATA_width, \
PWDATA_width=`PWDATA_width, \
PSTRB_width = `PSTRB_width, \
PADDR_width = `PADDT_width, \
PSELx_width = `PSELx_width \
)