`define PSELx_TIMEOUT_VAL 20
`define PSTRB_width 4
`define PWDATA_width 8 * `PSTRB_width
`define PRDATA_width  32
`define PADDR_width 32
`define PSELx_width 1
