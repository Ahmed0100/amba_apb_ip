`define IP_AMBA_APB_SLAVE_PARAM_DECL #(parameter PRDATA_width = `PRDATA_width, \
PRDATA_width=`PRDATA_width, \
PWDATA_width=`PWDATA_width, \
PSTRB_width = `PSTRB_width, \
PADDR_width = `PADDT_width, \
PSELx_width = `PSELx_width, \
WORD_LENGTH = `PRDATA_width, \
MEM_DEPTH = `MEM_ARRAY_SIZE_INT, \
APB_BASE_ADDR = `APB_base_addr \ 
)